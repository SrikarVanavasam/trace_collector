// pcie_ed_perf0.v

// Generated using ACDS version 24.3 212

`timescale 1 ps / 1 ps
module pcie_ed_perf0 (
		input  wire         coreclkout_hip,              //    coreclkout_hip.clk
		input  wire         p0_reset_status_n,           // p0_reset_status_n.reset_n
		input  wire         p1_reset_status_n,           // p1_reset_status_n.reset_n
		input  wire         p2_reset_status_n,           // p2_reset_status_n.reset_n
		input  wire         p3_reset_status_n,           // p3_reset_status_n.reset_n
		output wire         p0_rx_st_ready_o,            //         p0_rx_st0.ready
		input  wire [127:0] p0_rx_st0_data_i,            //                  .data
		input  wire         p0_rx_st0_sop_i,             //                  .startofpacket
		input  wire         p0_rx_st0_eop_i,             //                  .endofpacket
		input  wire         p0_rx_st0_dvalid_i,          //                  .valid
		input  wire [1:0]   p0_rx_st0_empty_i,           //                  .empty
		output wire         p1_rx_st_ready_o,            //         p1_rx_st0.ready
		input  wire [127:0] p1_rx_st0_data_i,            //                  .data
		input  wire         p1_rx_st0_sop_i,             //                  .startofpacket
		input  wire         p1_rx_st0_eop_i,             //                  .endofpacket
		input  wire         p1_rx_st0_dvalid_i,          //                  .valid
		input  wire [1:0]   p1_rx_st0_empty_i,           //                  .empty
		output wire         p2_rx_st_ready_o,            //         p2_rx_st0.ready
		input  wire [127:0] p2_rx_st0_data_i,            //                  .data
		input  wire         p2_rx_st0_sop_i,             //                  .startofpacket
		input  wire         p2_rx_st0_eop_i,             //                  .endofpacket
		input  wire         p2_rx_st0_dvalid_i,          //                  .valid
		input  wire [1:0]   p2_rx_st0_empty_i,           //                  .empty
		output wire         p3_rx_st_ready_o,            //         p3_rx_st0.ready
		input  wire [127:0] p3_rx_st0_data_i,            //                  .data
		input  wire         p3_rx_st0_sop_i,             //                  .startofpacket
		input  wire         p3_rx_st0_eop_i,             //                  .endofpacket
		input  wire         p3_rx_st0_dvalid_i,          //                  .valid
		input  wire [1:0]   p3_rx_st0_empty_i,           //                  .empty
		input  wire [127:0] p0_rx_st1_data_i,            //         p0_rx_st1.data
		input  wire         p0_rx_st1_sop_i,             //                  .startofpacket
		input  wire         p0_rx_st1_eop_i,             //                  .endofpacket
		input  wire         p0_rx_st1_dvalid_i,          //                  .valid
		input  wire [1:0]   p0_rx_st1_empty_i,           //                  .empty
		input  wire [127:0] p1_rx_st1_data_i,            //         p1_rx_st1.data
		input  wire         p1_rx_st1_sop_i,             //                  .startofpacket
		input  wire         p1_rx_st1_eop_i,             //                  .endofpacket
		input  wire         p1_rx_st1_dvalid_i,          //                  .valid
		input  wire [1:0]   p1_rx_st1_empty_i,           //                  .empty
		input  wire [127:0] p2_rx_st1_data_i,            //         p2_rx_st1.data
		input  wire         p2_rx_st1_sop_i,             //                  .startofpacket
		input  wire         p2_rx_st1_eop_i,             //                  .endofpacket
		input  wire         p2_rx_st1_dvalid_i,          //                  .valid
		input  wire [1:0]   p2_rx_st1_empty_i,           //                  .empty
		input  wire [127:0] p3_rx_st1_data_i,            //         p3_rx_st1.data
		input  wire         p3_rx_st1_sop_i,             //                  .startofpacket
		input  wire         p3_rx_st1_eop_i,             //                  .endofpacket
		input  wire         p3_rx_st1_dvalid_i,          //                  .valid
		input  wire [1:0]   p3_rx_st1_empty_i,           //                  .empty
		input  wire [127:0] p0_rx_st0_hdr_i,             //     p0_rx_st_misc.rx_st0_hdr
		input  wire [31:0]  p0_rx_st0_prefix_i,          //                  .rx_st0_prefix
		input  wire         p0_rx_st0_hvalid_i,          //                  .rx_st0_hvalid
		input  wire         p0_rx_st0_pvalid_i,          //                  .rx_st0_pvalid
		input  wire [2:0]   p0_rx_st0_bar_i,             //                  .rx_st0_bar
		input  wire [127:0] p0_rx_st1_hdr_i,             //                  .rx_st1_hdr
		input  wire [31:0]  p0_rx_st1_prefix_i,          //                  .rx_st1_prefix
		input  wire         p0_rx_st1_hvalid_i,          //                  .rx_st1_hvalid
		input  wire         p0_rx_st1_pvalid_i,          //                  .rx_st1_pvalid
		input  wire [2:0]   p0_rx_st1_bar_i,             //                  .rx_st1_bar
		output wire [2:0]   p0_rx_st_hcrdt_init_o,       //                  .rx_st_Hcrdt_init
		output wire [2:0]   p0_rx_st_hcrdt_update_o,     //                  .rx_st_Hcrdt_update
		output wire [5:0]   p0_rx_st_hcrdt_update_cnt_o, //                  .rx_st_Hcrdt_update_cnt
		input  wire [2:0]   p0_rx_st_hcrdt_init_ack_i,   //                  .rx_st_Hcrdt_init_ack
		output wire [2:0]   p0_rx_st_dcrdt_init_o,       //                  .rx_st_Dcrdt_init
		output wire [2:0]   p0_rx_st_dcrdt_update_o,     //                  .rx_st_Dcrdt_update
		output wire [11:0]  p0_rx_st_dcrdt_update_cnt_o, //                  .rx_st_Dcrdt_update_cnt
		input  wire [2:0]   p0_rx_st_dcrdt_init_ack_i,   //                  .rx_st_Dcrdt_init_ack
		input  wire [127:0] p1_rx_st0_hdr_i,             //     p1_rx_st_misc.rx_st0_hdr
		input  wire [31:0]  p1_rx_st0_prefix_i,          //                  .rx_st0_prefix
		input  wire         p1_rx_st0_hvalid_i,          //                  .rx_st0_hvalid
		input  wire         p1_rx_st0_pvalid_i,          //                  .rx_st0_pvalid
		input  wire [2:0]   p1_rx_st0_bar_i,             //                  .rx_st0_bar
		input  wire [127:0] p1_rx_st1_hdr_i,             //                  .rx_st1_hdr
		input  wire [31:0]  p1_rx_st1_prefix_i,          //                  .rx_st1_prefix
		input  wire         p1_rx_st1_hvalid_i,          //                  .rx_st1_hvalid
		input  wire         p1_rx_st1_pvalid_i,          //                  .rx_st1_pvalid
		input  wire [2:0]   p1_rx_st1_bar_i,             //                  .rx_st1_bar
		output wire [2:0]   p1_rx_st_hcrdt_init_o,       //                  .rx_st_Hcrdt_init
		output wire [2:0]   p1_rx_st_hcrdt_update_o,     //                  .rx_st_Hcrdt_update
		output wire [5:0]   p1_rx_st_hcrdt_update_cnt_o, //                  .rx_st_Hcrdt_update_cnt
		input  wire [2:0]   p1_rx_st_hcrdt_init_ack_i,   //                  .rx_st_Hcrdt_init_ack
		output wire [2:0]   p1_rx_st_dcrdt_init_o,       //                  .rx_st_Dcrdt_init
		output wire [2:0]   p1_rx_st_dcrdt_update_o,     //                  .rx_st_Dcrdt_update
		output wire [11:0]  p1_rx_st_dcrdt_update_cnt_o, //                  .rx_st_Dcrdt_update_cnt
		input  wire [2:0]   p1_rx_st_dcrdt_init_ack_i,   //                  .rx_st_Dcrdt_init_ack
		input  wire [127:0] p2_rx_st0_hdr_i,             //     p2_rx_st_misc.rx_st0_hdr
		input  wire [31:0]  p2_rx_st0_prefix_i,          //                  .rx_st0_prefix
		input  wire         p2_rx_st0_hvalid_i,          //                  .rx_st0_hvalid
		input  wire         p2_rx_st0_pvalid_i,          //                  .rx_st0_pvalid
		input  wire [2:0]   p2_rx_st0_bar_i,             //                  .rx_st0_bar
		input  wire [127:0] p2_rx_st1_hdr_i,             //                  .rx_st1_hdr
		input  wire [31:0]  p2_rx_st1_prefix_i,          //                  .rx_st1_prefix
		input  wire         p2_rx_st1_hvalid_i,          //                  .rx_st1_hvalid
		input  wire         p2_rx_st1_pvalid_i,          //                  .rx_st1_pvalid
		input  wire [2:0]   p2_rx_st1_bar_i,             //                  .rx_st1_bar
		output wire [2:0]   p2_rx_st_hcrdt_init_o,       //                  .rx_st_Hcrdt_init
		output wire [2:0]   p2_rx_st_hcrdt_update_o,     //                  .rx_st_Hcrdt_update
		output wire [5:0]   p2_rx_st_hcrdt_update_cnt_o, //                  .rx_st_Hcrdt_update_cnt
		input  wire [2:0]   p2_rx_st_hcrdt_init_ack_i,   //                  .rx_st_Hcrdt_init_ack
		output wire [2:0]   p2_rx_st_dcrdt_init_o,       //                  .rx_st_Dcrdt_init
		output wire [2:0]   p2_rx_st_dcrdt_update_o,     //                  .rx_st_Dcrdt_update
		output wire [11:0]  p2_rx_st_dcrdt_update_cnt_o, //                  .rx_st_Dcrdt_update_cnt
		input  wire [2:0]   p2_rx_st_dcrdt_init_ack_i,   //                  .rx_st_Dcrdt_init_ack
		input  wire [127:0] p3_rx_st0_hdr_i,             //     p3_rx_st_misc.rx_st0_hdr
		input  wire [31:0]  p3_rx_st0_prefix_i,          //                  .rx_st0_prefix
		input  wire         p3_rx_st0_hvalid_i,          //                  .rx_st0_hvalid
		input  wire         p3_rx_st0_pvalid_i,          //                  .rx_st0_pvalid
		input  wire [2:0]   p3_rx_st0_bar_i,             //                  .rx_st0_bar
		input  wire [127:0] p3_rx_st1_hdr_i,             //                  .rx_st1_hdr
		input  wire [31:0]  p3_rx_st1_prefix_i,          //                  .rx_st1_prefix
		input  wire         p3_rx_st1_hvalid_i,          //                  .rx_st1_hvalid
		input  wire         p3_rx_st1_pvalid_i,          //                  .rx_st1_pvalid
		input  wire [2:0]   p3_rx_st1_bar_i,             //                  .rx_st1_bar
		output wire [2:0]   p3_rx_st_hcrdt_init_o,       //                  .rx_st_Hcrdt_init
		output wire [2:0]   p3_rx_st_hcrdt_update_o,     //                  .rx_st_Hcrdt_update
		output wire [5:0]   p3_rx_st_hcrdt_update_cnt_o, //                  .rx_st_Hcrdt_update_cnt
		input  wire [2:0]   p3_rx_st_hcrdt_init_ack_i,   //                  .rx_st_Hcrdt_init_ack
		output wire [2:0]   p3_rx_st_dcrdt_init_o,       //                  .rx_st_Dcrdt_init
		output wire [2:0]   p3_rx_st_dcrdt_update_o,     //                  .rx_st_Dcrdt_update
		output wire [11:0]  p3_rx_st_dcrdt_update_cnt_o, //                  .rx_st_Dcrdt_update_cnt
		input  wire [2:0]   p3_rx_st_dcrdt_init_ack_i,   //                  .rx_st_Dcrdt_init_ack
		input  wire [2:0]   p0_tx_st_hcrdt_init_i,       //     p0_tx_st_misc.tx_st_Hcrdt_init
		input  wire [2:0]   p0_tx_st_hcrdt_update_i,     //                  .tx_st_Hcrdt_update
		input  wire [5:0]   p0_tx_st_hcrdt_update_cnt_i, //                  .tx_st_Hcrdt_update_cnt
		output wire [2:0]   p0_tx_st_hcrdt_init_ack_o,   //                  .tx_st_Hcrdtt_init_ack
		input  wire [2:0]   p0_tx_st_dcrdt_init_i,       //                  .tx_st_Dcrdt_init
		input  wire [2:0]   p0_tx_st_dcrdt_update_i,     //                  .tx_st_Dcrdt_update
		input  wire [11:0]  p0_tx_st_dcrdt_update_cnt_i, //                  .tx_st_Dcrdt_update_cnt
		output wire [2:0]   p0_tx_st_dcrdt_init_ack_o,   //                  .tx_st_Dcrdt_init_ack
		output wire [127:0] p0_tx_st0_hdr_o,             //                  .tx_st0_hdr
		output wire [31:0]  p0_tx_st0_prefix_o,          //                  .tx_st0_prefix
		output wire         p0_tx_st0_hvalid_o,          //                  .tx_st0_hvalid
		output wire         p0_tx_st0_pvalid_o,          //                  .tx_st0_pvalid
		output wire [127:0] p0_tx_st1_hdr_o,             //                  .tx_st1_hdr
		output wire [31:0]  p0_tx_st1_prefix_o,          //                  .tx_st1_prefix
		output wire         p0_tx_st1_hvalid_o,          //                  .tx_st1_hvalid
		output wire         p0_tx_st1_pvalid_o,          //                  .tx_st1_pvalid
		input  wire [2:0]   p1_tx_st_hcrdt_init_i,       //     p1_tx_st_misc.tx_st_Hcrdt_init
		input  wire [2:0]   p1_tx_st_hcrdt_update_i,     //                  .tx_st_Hcrdt_update
		input  wire [5:0]   p1_tx_st_hcrdt_update_cnt_i, //                  .tx_st_Hcrdt_update_cnt
		output wire [2:0]   p1_tx_st_hcrdt_init_ack_o,   //                  .tx_st_Hcrdtt_init_ack
		input  wire [2:0]   p1_tx_st_dcrdt_init_i,       //                  .tx_st_Dcrdt_init
		input  wire [2:0]   p1_tx_st_dcrdt_update_i,     //                  .tx_st_Dcrdt_update
		input  wire [11:0]  p1_tx_st_dcrdt_update_cnt_i, //                  .tx_st_Dcrdt_update_cnt
		output wire [2:0]   p1_tx_st_dcrdt_init_ack_o,   //                  .tx_st_Dcrdt_init_ack
		output wire [127:0] p1_tx_st0_hdr_o,             //                  .tx_st0_hdr
		output wire [31:0]  p1_tx_st0_prefix_o,          //                  .tx_st0_prefix
		output wire         p1_tx_st0_hvalid_o,          //                  .tx_st0_hvalid
		output wire         p1_tx_st0_pvalid_o,          //                  .tx_st0_pvalid
		output wire [127:0] p1_tx_st1_hdr_o,             //                  .tx_st1_hdr
		output wire [31:0]  p1_tx_st1_prefix_o,          //                  .tx_st1_prefix
		output wire         p1_tx_st1_hvalid_o,          //                  .tx_st1_hvalid
		output wire         p1_tx_st1_pvalid_o,          //                  .tx_st1_pvalid
		input  wire [2:0]   p2_tx_st_hcrdt_init_i,       //     p2_tx_st_misc.tx_st_Hcrdt_init
		input  wire [2:0]   p2_tx_st_hcrdt_update_i,     //                  .tx_st_Hcrdt_update
		input  wire [5:0]   p2_tx_st_hcrdt_update_cnt_i, //                  .tx_st_Hcrdt_update_cnt
		output wire [2:0]   p2_tx_st_hcrdt_init_ack_o,   //                  .tx_st_Hcrdtt_init_ack
		input  wire [2:0]   p2_tx_st_dcrdt_init_i,       //                  .tx_st_Dcrdt_init
		input  wire [2:0]   p2_tx_st_dcrdt_update_i,     //                  .tx_st_Dcrdt_update
		input  wire [11:0]  p2_tx_st_dcrdt_update_cnt_i, //                  .tx_st_Dcrdt_update_cnt
		output wire [2:0]   p2_tx_st_dcrdt_init_ack_o,   //                  .tx_st_Dcrdt_init_ack
		output wire [127:0] p2_tx_st0_hdr_o,             //                  .tx_st0_hdr
		output wire [31:0]  p2_tx_st0_prefix_o,          //                  .tx_st0_prefix
		output wire         p2_tx_st0_hvalid_o,          //                  .tx_st0_hvalid
		output wire         p2_tx_st0_pvalid_o,          //                  .tx_st0_pvalid
		output wire [127:0] p2_tx_st1_hdr_o,             //                  .tx_st1_hdr
		output wire [31:0]  p2_tx_st1_prefix_o,          //                  .tx_st1_prefix
		output wire         p2_tx_st1_hvalid_o,          //                  .tx_st1_hvalid
		output wire         p2_tx_st1_pvalid_o,          //                  .tx_st1_pvalid
		input  wire [2:0]   p3_tx_st_hcrdt_init_i,       //     p3_tx_st_misc.tx_st_Hcrdt_init
		input  wire [2:0]   p3_tx_st_hcrdt_update_i,     //                  .tx_st_Hcrdt_update
		input  wire [5:0]   p3_tx_st_hcrdt_update_cnt_i, //                  .tx_st_Hcrdt_update_cnt
		output wire [2:0]   p3_tx_st_hcrdt_init_ack_o,   //                  .tx_st_Hcrdtt_init_ack
		input  wire [2:0]   p3_tx_st_dcrdt_init_i,       //                  .tx_st_Dcrdt_init
		input  wire [2:0]   p3_tx_st_dcrdt_update_i,     //                  .tx_st_Dcrdt_update
		input  wire [11:0]  p3_tx_st_dcrdt_update_cnt_i, //                  .tx_st_Dcrdt_update_cnt
		output wire [2:0]   p3_tx_st_dcrdt_init_ack_o,   //                  .tx_st_Dcrdt_init_ack
		output wire [127:0] p3_tx_st0_hdr_o,             //                  .tx_st0_hdr
		output wire [31:0]  p3_tx_st0_prefix_o,          //                  .tx_st0_prefix
		output wire         p3_tx_st0_hvalid_o,          //                  .tx_st0_hvalid
		output wire         p3_tx_st0_pvalid_o,          //                  .tx_st0_pvalid
		output wire [127:0] p3_tx_st1_hdr_o,             //                  .tx_st1_hdr
		output wire [31:0]  p3_tx_st1_prefix_o,          //                  .tx_st1_prefix
		output wire         p3_tx_st1_hvalid_o,          //                  .tx_st1_hvalid
		output wire         p3_tx_st1_pvalid_o,          //                  .tx_st1_pvalid
		input  wire         p0_tx_st0_ready_i,           //         p0_tx_st0.ready
		output wire [127:0] p0_tx_st0_data_o,            //                  .data
		output wire         p0_tx_st0_sop_o,             //                  .startofpacket
		output wire         p0_tx_st0_eop_o,             //                  .endofpacket
		output wire         p0_tx_st0_dvalid_o,          //                  .valid
		input  wire         p1_tx_st0_ready_i,           //         p1_tx_st0.ready
		output wire [127:0] p1_tx_st0_data_o,            //                  .data
		output wire         p1_tx_st0_sop_o,             //                  .startofpacket
		output wire         p1_tx_st0_eop_o,             //                  .endofpacket
		output wire         p1_tx_st0_dvalid_o,          //                  .valid
		input  wire         p2_tx_st0_ready_i,           //         p2_tx_st0.ready
		output wire [127:0] p2_tx_st0_data_o,            //                  .data
		output wire         p2_tx_st0_sop_o,             //                  .startofpacket
		output wire         p2_tx_st0_eop_o,             //                  .endofpacket
		output wire         p2_tx_st0_dvalid_o,          //                  .valid
		input  wire         p3_tx_st0_ready_i,           //         p3_tx_st0.ready
		output wire [127:0] p3_tx_st0_data_o,            //                  .data
		output wire         p3_tx_st0_sop_o,             //                  .startofpacket
		output wire         p3_tx_st0_eop_o,             //                  .endofpacket
		output wire         p3_tx_st0_dvalid_o,          //                  .valid
		output wire [127:0] p0_tx_st1_data_o,            //         p0_tx_st1.data
		output wire         p0_tx_st1_sop_o,             //                  .startofpacket
		output wire         p0_tx_st1_eop_o,             //                  .endofpacket
		output wire         p0_tx_st1_dvalid_o,          //                  .valid
		output wire [127:0] p1_tx_st1_data_o,            //         p1_tx_st1.data
		output wire         p1_tx_st1_sop_o,             //                  .startofpacket
		output wire         p1_tx_st1_eop_o,             //                  .endofpacket
		output wire         p1_tx_st1_dvalid_o,          //                  .valid
		output wire [127:0] p2_tx_st1_data_o,            //         p2_tx_st1.data
		output wire         p2_tx_st1_sop_o,             //                  .startofpacket
		output wire         p2_tx_st1_eop_o,             //                  .endofpacket
		output wire         p2_tx_st1_dvalid_o,          //                  .valid
		output wire [127:0] p3_tx_st1_data_o,            //         p3_tx_st1.data
		output wire         p3_tx_st1_sop_o,             //                  .startofpacket
		output wire         p3_tx_st1_eop_o,             //                  .endofpacket
		output wire         p3_tx_st1_dvalid_o,          //                  .valid

    // Between CXL and PCIe
    input logic                         trace_valid_0,
    input logic                         trace_valid_1,
    input logic [511:0]                 trace_data_0,
    input logic [511:0]                 trace_data_1,
    input logic [63:0]                  trace_buffer_base_addr_0,
    input logic [63:0]                  trace_buffer_base_addr_1,
    input logic [63:0]                  trace_buffer_size_0,
    input logic [63:0]                  trace_buffer_size_1,
    input logic [63:0]                  control_register_0,
    input logic [63:0]                  control_register_1,
    output  logic [63:0]                  dropped_traces_0,
    output  logic [63:0]                  dropped_traces_1,
    output  logic [63:0]                  written_traces_0,
    output  logic [63:0]                  written_traces_1
	);

	intel_pcie_perf_ed_gen5 #(
		.LANE_MODE ("PCIE_X4X4")
	) perf0 (
		.coreclkout_hip              (coreclkout_hip),              //   input,    width = 1,    coreclkout_hip.clk
		.p0_reset_status_n           (p0_reset_status_n),           //   input,    width = 1, p0_reset_status_n.reset_n
		.p1_reset_status_n           (p1_reset_status_n),           //   input,    width = 1, p1_reset_status_n.reset_n
		.p2_reset_status_n           (p2_reset_status_n),           //   input,    width = 1, p2_reset_status_n.reset_n
		.p3_reset_status_n           (p3_reset_status_n),           //   input,    width = 1, p3_reset_status_n.reset_n
		.p0_rx_st_ready_o            (p0_rx_st_ready_o),            //  output,    width = 1,         p0_rx_st0.ready
		.p0_rx_st0_data_i            (p0_rx_st0_data_i),            //   input,  width = 128,                  .data
		.p0_rx_st0_sop_i             (p0_rx_st0_sop_i),             //   input,    width = 1,                  .startofpacket
		.p0_rx_st0_eop_i             (p0_rx_st0_eop_i),             //   input,    width = 1,                  .endofpacket
		.p0_rx_st0_dvalid_i          (p0_rx_st0_dvalid_i),          //   input,    width = 1,                  .valid
		.p0_rx_st0_empty_i           (p0_rx_st0_empty_i),           //   input,    width = 2,                  .empty
		.p1_rx_st_ready_o            (p1_rx_st_ready_o),            //  output,    width = 1,         p1_rx_st0.ready
		.p1_rx_st0_data_i            (p1_rx_st0_data_i),            //   input,  width = 128,                  .data
		.p1_rx_st0_sop_i             (p1_rx_st0_sop_i),             //   input,    width = 1,                  .startofpacket
		.p1_rx_st0_eop_i             (p1_rx_st0_eop_i),             //   input,    width = 1,                  .endofpacket
		.p1_rx_st0_dvalid_i          (p1_rx_st0_dvalid_i),          //   input,    width = 1,                  .valid
		.p1_rx_st0_empty_i           (p1_rx_st0_empty_i),           //   input,    width = 2,                  .empty
		.p2_rx_st_ready_o            (p2_rx_st_ready_o),            //  output,    width = 1,         p2_rx_st0.ready
		.p2_rx_st0_data_i            (p2_rx_st0_data_i),            //   input,  width = 128,                  .data
		.p2_rx_st0_sop_i             (p2_rx_st0_sop_i),             //   input,    width = 1,                  .startofpacket
		.p2_rx_st0_eop_i             (p2_rx_st0_eop_i),             //   input,    width = 1,                  .endofpacket
		.p2_rx_st0_dvalid_i          (p2_rx_st0_dvalid_i),          //   input,    width = 1,                  .valid
		.p2_rx_st0_empty_i           (p2_rx_st0_empty_i),           //   input,    width = 2,                  .empty
		.p3_rx_st_ready_o            (p3_rx_st_ready_o),            //  output,    width = 1,         p3_rx_st0.ready
		.p3_rx_st0_data_i            (p3_rx_st0_data_i),            //   input,  width = 128,                  .data
		.p3_rx_st0_sop_i             (p3_rx_st0_sop_i),             //   input,    width = 1,                  .startofpacket
		.p3_rx_st0_eop_i             (p3_rx_st0_eop_i),             //   input,    width = 1,                  .endofpacket
		.p3_rx_st0_dvalid_i          (p3_rx_st0_dvalid_i),          //   input,    width = 1,                  .valid
		.p3_rx_st0_empty_i           (p3_rx_st0_empty_i),           //   input,    width = 2,                  .empty
		.p0_rx_st1_data_i            (p0_rx_st1_data_i),            //   input,  width = 128,         p0_rx_st1.data
		.p0_rx_st1_sop_i             (p0_rx_st1_sop_i),             //   input,    width = 1,                  .startofpacket
		.p0_rx_st1_eop_i             (p0_rx_st1_eop_i),             //   input,    width = 1,                  .endofpacket
		.p0_rx_st1_dvalid_i          (p0_rx_st1_dvalid_i),          //   input,    width = 1,                  .valid
		.p0_rx_st1_empty_i           (p0_rx_st1_empty_i),           //   input,    width = 2,                  .empty
		.p1_rx_st1_data_i            (p1_rx_st1_data_i),            //   input,  width = 128,         p1_rx_st1.data
		.p1_rx_st1_sop_i             (p1_rx_st1_sop_i),             //   input,    width = 1,                  .startofpacket
		.p1_rx_st1_eop_i             (p1_rx_st1_eop_i),             //   input,    width = 1,                  .endofpacket
		.p1_rx_st1_dvalid_i          (p1_rx_st1_dvalid_i),          //   input,    width = 1,                  .valid
		.p1_rx_st1_empty_i           (p1_rx_st1_empty_i),           //   input,    width = 2,                  .empty
		.p2_rx_st1_data_i            (p2_rx_st1_data_i),            //   input,  width = 128,         p2_rx_st1.data
		.p2_rx_st1_sop_i             (p2_rx_st1_sop_i),             //   input,    width = 1,                  .startofpacket
		.p2_rx_st1_eop_i             (p2_rx_st1_eop_i),             //   input,    width = 1,                  .endofpacket
		.p2_rx_st1_dvalid_i          (p2_rx_st1_dvalid_i),          //   input,    width = 1,                  .valid
		.p2_rx_st1_empty_i           (p2_rx_st1_empty_i),           //   input,    width = 2,                  .empty
		.p3_rx_st1_data_i            (p3_rx_st1_data_i),            //   input,  width = 128,         p3_rx_st1.data
		.p3_rx_st1_sop_i             (p3_rx_st1_sop_i),             //   input,    width = 1,                  .startofpacket
		.p3_rx_st1_eop_i             (p3_rx_st1_eop_i),             //   input,    width = 1,                  .endofpacket
		.p3_rx_st1_dvalid_i          (p3_rx_st1_dvalid_i),          //   input,    width = 1,                  .valid
		.p3_rx_st1_empty_i           (p3_rx_st1_empty_i),           //   input,    width = 2,                  .empty
		.p0_rx_st0_hdr_i             (p0_rx_st0_hdr_i),             //   input,  width = 128,     p0_rx_st_misc.rx_st0_hdr
		.p0_rx_st0_prefix_i          (p0_rx_st0_prefix_i),          //   input,   width = 32,                  .rx_st0_prefix
		.p0_rx_st0_hvalid_i          (p0_rx_st0_hvalid_i),          //   input,    width = 1,                  .rx_st0_hvalid
		.p0_rx_st0_pvalid_i          (p0_rx_st0_pvalid_i),          //   input,    width = 1,                  .rx_st0_pvalid
		.p0_rx_st0_bar_i             (p0_rx_st0_bar_i),             //   input,    width = 3,                  .rx_st0_bar
		.p0_rx_st1_hdr_i             (p0_rx_st1_hdr_i),             //   input,  width = 128,                  .rx_st1_hdr
		.p0_rx_st1_prefix_i          (p0_rx_st1_prefix_i),          //   input,   width = 32,                  .rx_st1_prefix
		.p0_rx_st1_hvalid_i          (p0_rx_st1_hvalid_i),          //   input,    width = 1,                  .rx_st1_hvalid
		.p0_rx_st1_pvalid_i          (p0_rx_st1_pvalid_i),          //   input,    width = 1,                  .rx_st1_pvalid
		.p0_rx_st1_bar_i             (p0_rx_st1_bar_i),             //   input,    width = 3,                  .rx_st1_bar
		.p0_rx_st_hcrdt_init_o       (p0_rx_st_hcrdt_init_o),       //  output,    width = 3,                  .rx_st_Hcrdt_init
		.p0_rx_st_hcrdt_update_o     (p0_rx_st_hcrdt_update_o),     //  output,    width = 3,                  .rx_st_Hcrdt_update
		.p0_rx_st_hcrdt_update_cnt_o (p0_rx_st_hcrdt_update_cnt_o), //  output,    width = 6,                  .rx_st_Hcrdt_update_cnt
		.p0_rx_st_hcrdt_init_ack_i   (p0_rx_st_hcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Hcrdt_init_ack
		.p0_rx_st_dcrdt_init_o       (p0_rx_st_dcrdt_init_o),       //  output,    width = 3,                  .rx_st_Dcrdt_init
		.p0_rx_st_dcrdt_update_o     (p0_rx_st_dcrdt_update_o),     //  output,    width = 3,                  .rx_st_Dcrdt_update
		.p0_rx_st_dcrdt_update_cnt_o (p0_rx_st_dcrdt_update_cnt_o), //  output,   width = 12,                  .rx_st_Dcrdt_update_cnt
		.p0_rx_st_dcrdt_init_ack_i   (p0_rx_st_dcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Dcrdt_init_ack
		.p1_rx_st0_hdr_i             (p1_rx_st0_hdr_i),             //   input,  width = 128,     p1_rx_st_misc.rx_st0_hdr
		.p1_rx_st0_prefix_i          (p1_rx_st0_prefix_i),          //   input,   width = 32,                  .rx_st0_prefix
		.p1_rx_st0_hvalid_i          (p1_rx_st0_hvalid_i),          //   input,    width = 1,                  .rx_st0_hvalid
		.p1_rx_st0_pvalid_i          (p1_rx_st0_pvalid_i),          //   input,    width = 1,                  .rx_st0_pvalid
		.p1_rx_st0_bar_i             (p1_rx_st0_bar_i),             //   input,    width = 3,                  .rx_st0_bar
		.p1_rx_st1_hdr_i             (p1_rx_st1_hdr_i),             //   input,  width = 128,                  .rx_st1_hdr
		.p1_rx_st1_prefix_i          (p1_rx_st1_prefix_i),          //   input,   width = 32,                  .rx_st1_prefix
		.p1_rx_st1_hvalid_i          (p1_rx_st1_hvalid_i),          //   input,    width = 1,                  .rx_st1_hvalid
		.p1_rx_st1_pvalid_i          (p1_rx_st1_pvalid_i),          //   input,    width = 1,                  .rx_st1_pvalid
		.p1_rx_st1_bar_i             (p1_rx_st1_bar_i),             //   input,    width = 3,                  .rx_st1_bar
		.p1_rx_st_hcrdt_init_o       (p1_rx_st_hcrdt_init_o),       //  output,    width = 3,                  .rx_st_Hcrdt_init
		.p1_rx_st_hcrdt_update_o     (p1_rx_st_hcrdt_update_o),     //  output,    width = 3,                  .rx_st_Hcrdt_update
		.p1_rx_st_hcrdt_update_cnt_o (p1_rx_st_hcrdt_update_cnt_o), //  output,    width = 6,                  .rx_st_Hcrdt_update_cnt
		.p1_rx_st_hcrdt_init_ack_i   (p1_rx_st_hcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Hcrdt_init_ack
		.p1_rx_st_dcrdt_init_o       (p1_rx_st_dcrdt_init_o),       //  output,    width = 3,                  .rx_st_Dcrdt_init
		.p1_rx_st_dcrdt_update_o     (p1_rx_st_dcrdt_update_o),     //  output,    width = 3,                  .rx_st_Dcrdt_update
		.p1_rx_st_dcrdt_update_cnt_o (p1_rx_st_dcrdt_update_cnt_o), //  output,   width = 12,                  .rx_st_Dcrdt_update_cnt
		.p1_rx_st_dcrdt_init_ack_i   (p1_rx_st_dcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Dcrdt_init_ack
		.p2_rx_st0_hdr_i             (p2_rx_st0_hdr_i),             //   input,  width = 128,     p2_rx_st_misc.rx_st0_hdr
		.p2_rx_st0_prefix_i          (p2_rx_st0_prefix_i),          //   input,   width = 32,                  .rx_st0_prefix
		.p2_rx_st0_hvalid_i          (p2_rx_st0_hvalid_i),          //   input,    width = 1,                  .rx_st0_hvalid
		.p2_rx_st0_pvalid_i          (p2_rx_st0_pvalid_i),          //   input,    width = 1,                  .rx_st0_pvalid
		.p2_rx_st0_bar_i             (p2_rx_st0_bar_i),             //   input,    width = 3,                  .rx_st0_bar
		.p2_rx_st1_hdr_i             (p2_rx_st1_hdr_i),             //   input,  width = 128,                  .rx_st1_hdr
		.p2_rx_st1_prefix_i          (p2_rx_st1_prefix_i),          //   input,   width = 32,                  .rx_st1_prefix
		.p2_rx_st1_hvalid_i          (p2_rx_st1_hvalid_i),          //   input,    width = 1,                  .rx_st1_hvalid
		.p2_rx_st1_pvalid_i          (p2_rx_st1_pvalid_i),          //   input,    width = 1,                  .rx_st1_pvalid
		.p2_rx_st1_bar_i             (p2_rx_st1_bar_i),             //   input,    width = 3,                  .rx_st1_bar
		.p2_rx_st_hcrdt_init_o       (p2_rx_st_hcrdt_init_o),       //  output,    width = 3,                  .rx_st_Hcrdt_init
		.p2_rx_st_hcrdt_update_o     (p2_rx_st_hcrdt_update_o),     //  output,    width = 3,                  .rx_st_Hcrdt_update
		.p2_rx_st_hcrdt_update_cnt_o (p2_rx_st_hcrdt_update_cnt_o), //  output,    width = 6,                  .rx_st_Hcrdt_update_cnt
		.p2_rx_st_hcrdt_init_ack_i   (p2_rx_st_hcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Hcrdt_init_ack
		.p2_rx_st_dcrdt_init_o       (p2_rx_st_dcrdt_init_o),       //  output,    width = 3,                  .rx_st_Dcrdt_init
		.p2_rx_st_dcrdt_update_o     (p2_rx_st_dcrdt_update_o),     //  output,    width = 3,                  .rx_st_Dcrdt_update
		.p2_rx_st_dcrdt_update_cnt_o (p2_rx_st_dcrdt_update_cnt_o), //  output,   width = 12,                  .rx_st_Dcrdt_update_cnt
		.p2_rx_st_dcrdt_init_ack_i   (p2_rx_st_dcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Dcrdt_init_ack
		.p3_rx_st0_hdr_i             (p3_rx_st0_hdr_i),             //   input,  width = 128,     p3_rx_st_misc.rx_st0_hdr
		.p3_rx_st0_prefix_i          (p3_rx_st0_prefix_i),          //   input,   width = 32,                  .rx_st0_prefix
		.p3_rx_st0_hvalid_i          (p3_rx_st0_hvalid_i),          //   input,    width = 1,                  .rx_st0_hvalid
		.p3_rx_st0_pvalid_i          (p3_rx_st0_pvalid_i),          //   input,    width = 1,                  .rx_st0_pvalid
		.p3_rx_st0_bar_i             (p3_rx_st0_bar_i),             //   input,    width = 3,                  .rx_st0_bar
		.p3_rx_st1_hdr_i             (p3_rx_st1_hdr_i),             //   input,  width = 128,                  .rx_st1_hdr
		.p3_rx_st1_prefix_i          (p3_rx_st1_prefix_i),          //   input,   width = 32,                  .rx_st1_prefix
		.p3_rx_st1_hvalid_i          (p3_rx_st1_hvalid_i),          //   input,    width = 1,                  .rx_st1_hvalid
		.p3_rx_st1_pvalid_i          (p3_rx_st1_pvalid_i),          //   input,    width = 1,                  .rx_st1_pvalid
		.p3_rx_st1_bar_i             (p3_rx_st1_bar_i),             //   input,    width = 3,                  .rx_st1_bar
		.p3_rx_st_hcrdt_init_o       (p3_rx_st_hcrdt_init_o),       //  output,    width = 3,                  .rx_st_Hcrdt_init
		.p3_rx_st_hcrdt_update_o     (p3_rx_st_hcrdt_update_o),     //  output,    width = 3,                  .rx_st_Hcrdt_update
		.p3_rx_st_hcrdt_update_cnt_o (p3_rx_st_hcrdt_update_cnt_o), //  output,    width = 6,                  .rx_st_Hcrdt_update_cnt
		.p3_rx_st_hcrdt_init_ack_i   (p3_rx_st_hcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Hcrdt_init_ack
		.p3_rx_st_dcrdt_init_o       (p3_rx_st_dcrdt_init_o),       //  output,    width = 3,                  .rx_st_Dcrdt_init
		.p3_rx_st_dcrdt_update_o     (p3_rx_st_dcrdt_update_o),     //  output,    width = 3,                  .rx_st_Dcrdt_update
		.p3_rx_st_dcrdt_update_cnt_o (p3_rx_st_dcrdt_update_cnt_o), //  output,   width = 12,                  .rx_st_Dcrdt_update_cnt
		.p3_rx_st_dcrdt_init_ack_i   (p3_rx_st_dcrdt_init_ack_i),   //   input,    width = 3,                  .rx_st_Dcrdt_init_ack
		.p0_tx_st_hcrdt_init_i       (p0_tx_st_hcrdt_init_i),       //   input,    width = 3,     p0_tx_st_misc.tx_st_Hcrdt_init
		.p0_tx_st_hcrdt_update_i     (p0_tx_st_hcrdt_update_i),     //   input,    width = 3,                  .tx_st_Hcrdt_update
		.p0_tx_st_hcrdt_update_cnt_i (p0_tx_st_hcrdt_update_cnt_i), //   input,    width = 6,                  .tx_st_Hcrdt_update_cnt
		.p0_tx_st_hcrdt_init_ack_o   (p0_tx_st_hcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Hcrdtt_init_ack
		.p0_tx_st_dcrdt_init_i       (p0_tx_st_dcrdt_init_i),       //   input,    width = 3,                  .tx_st_Dcrdt_init
		.p0_tx_st_dcrdt_update_i     (p0_tx_st_dcrdt_update_i),     //   input,    width = 3,                  .tx_st_Dcrdt_update
		.p0_tx_st_dcrdt_update_cnt_i (p0_tx_st_dcrdt_update_cnt_i), //   input,   width = 12,                  .tx_st_Dcrdt_update_cnt
		.p0_tx_st_dcrdt_init_ack_o   (p0_tx_st_dcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Dcrdt_init_ack
		.p0_tx_st0_hdr_o             (p0_tx_st0_hdr_o),             //  output,  width = 128,                  .tx_st0_hdr
		.p0_tx_st0_prefix_o          (p0_tx_st0_prefix_o),          //  output,   width = 32,                  .tx_st0_prefix
		.p0_tx_st0_hvalid_o          (p0_tx_st0_hvalid_o),          //  output,    width = 1,                  .tx_st0_hvalid
		.p0_tx_st0_pvalid_o          (p0_tx_st0_pvalid_o),          //  output,    width = 1,                  .tx_st0_pvalid
		.p0_tx_st1_hdr_o             (p0_tx_st1_hdr_o),             //  output,  width = 128,                  .tx_st1_hdr
		.p0_tx_st1_prefix_o          (p0_tx_st1_prefix_o),          //  output,   width = 32,                  .tx_st1_prefix
		.p0_tx_st1_hvalid_o          (p0_tx_st1_hvalid_o),          //  output,    width = 1,                  .tx_st1_hvalid
		.p0_tx_st1_pvalid_o          (p0_tx_st1_pvalid_o),          //  output,    width = 1,                  .tx_st1_pvalid
		.p1_tx_st_hcrdt_init_i       (p1_tx_st_hcrdt_init_i),       //   input,    width = 3,     p1_tx_st_misc.tx_st_Hcrdt_init
		.p1_tx_st_hcrdt_update_i     (p1_tx_st_hcrdt_update_i),     //   input,    width = 3,                  .tx_st_Hcrdt_update
		.p1_tx_st_hcrdt_update_cnt_i (p1_tx_st_hcrdt_update_cnt_i), //   input,    width = 6,                  .tx_st_Hcrdt_update_cnt
		.p1_tx_st_hcrdt_init_ack_o   (p1_tx_st_hcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Hcrdtt_init_ack
		.p1_tx_st_dcrdt_init_i       (p1_tx_st_dcrdt_init_i),       //   input,    width = 3,                  .tx_st_Dcrdt_init
		.p1_tx_st_dcrdt_update_i     (p1_tx_st_dcrdt_update_i),     //   input,    width = 3,                  .tx_st_Dcrdt_update
		.p1_tx_st_dcrdt_update_cnt_i (p1_tx_st_dcrdt_update_cnt_i), //   input,   width = 12,                  .tx_st_Dcrdt_update_cnt
		.p1_tx_st_dcrdt_init_ack_o   (p1_tx_st_dcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Dcrdt_init_ack
		.p1_tx_st0_hdr_o             (p1_tx_st0_hdr_o),             //  output,  width = 128,                  .tx_st0_hdr
		.p1_tx_st0_prefix_o          (p1_tx_st0_prefix_o),          //  output,   width = 32,                  .tx_st0_prefix
		.p1_tx_st0_hvalid_o          (p1_tx_st0_hvalid_o),          //  output,    width = 1,                  .tx_st0_hvalid
		.p1_tx_st0_pvalid_o          (p1_tx_st0_pvalid_o),          //  output,    width = 1,                  .tx_st0_pvalid
		.p1_tx_st1_hdr_o             (p1_tx_st1_hdr_o),             //  output,  width = 128,                  .tx_st1_hdr
		.p1_tx_st1_prefix_o          (p1_tx_st1_prefix_o),          //  output,   width = 32,                  .tx_st1_prefix
		.p1_tx_st1_hvalid_o          (p1_tx_st1_hvalid_o),          //  output,    width = 1,                  .tx_st1_hvalid
		.p1_tx_st1_pvalid_o          (p1_tx_st1_pvalid_o),          //  output,    width = 1,                  .tx_st1_pvalid
		.p2_tx_st_hcrdt_init_i       (p2_tx_st_hcrdt_init_i),       //   input,    width = 3,     p2_tx_st_misc.tx_st_Hcrdt_init
		.p2_tx_st_hcrdt_update_i     (p2_tx_st_hcrdt_update_i),     //   input,    width = 3,                  .tx_st_Hcrdt_update
		.p2_tx_st_hcrdt_update_cnt_i (p2_tx_st_hcrdt_update_cnt_i), //   input,    width = 6,                  .tx_st_Hcrdt_update_cnt
		.p2_tx_st_hcrdt_init_ack_o   (p2_tx_st_hcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Hcrdtt_init_ack
		.p2_tx_st_dcrdt_init_i       (p2_tx_st_dcrdt_init_i),       //   input,    width = 3,                  .tx_st_Dcrdt_init
		.p2_tx_st_dcrdt_update_i     (p2_tx_st_dcrdt_update_i),     //   input,    width = 3,                  .tx_st_Dcrdt_update
		.p2_tx_st_dcrdt_update_cnt_i (p2_tx_st_dcrdt_update_cnt_i), //   input,   width = 12,                  .tx_st_Dcrdt_update_cnt
		.p2_tx_st_dcrdt_init_ack_o   (p2_tx_st_dcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Dcrdt_init_ack
		.p2_tx_st0_hdr_o             (p2_tx_st0_hdr_o),             //  output,  width = 128,                  .tx_st0_hdr
		.p2_tx_st0_prefix_o          (p2_tx_st0_prefix_o),          //  output,   width = 32,                  .tx_st0_prefix
		.p2_tx_st0_hvalid_o          (p2_tx_st0_hvalid_o),          //  output,    width = 1,                  .tx_st0_hvalid
		.p2_tx_st0_pvalid_o          (p2_tx_st0_pvalid_o),          //  output,    width = 1,                  .tx_st0_pvalid
		.p2_tx_st1_hdr_o             (p2_tx_st1_hdr_o),             //  output,  width = 128,                  .tx_st1_hdr
		.p2_tx_st1_prefix_o          (p2_tx_st1_prefix_o),          //  output,   width = 32,                  .tx_st1_prefix
		.p2_tx_st1_hvalid_o          (p2_tx_st1_hvalid_o),          //  output,    width = 1,                  .tx_st1_hvalid
		.p2_tx_st1_pvalid_o          (p2_tx_st1_pvalid_o),          //  output,    width = 1,                  .tx_st1_pvalid
		.p3_tx_st_hcrdt_init_i       (p3_tx_st_hcrdt_init_i),       //   input,    width = 3,     p3_tx_st_misc.tx_st_Hcrdt_init
		.p3_tx_st_hcrdt_update_i     (p3_tx_st_hcrdt_update_i),     //   input,    width = 3,                  .tx_st_Hcrdt_update
		.p3_tx_st_hcrdt_update_cnt_i (p3_tx_st_hcrdt_update_cnt_i), //   input,    width = 6,                  .tx_st_Hcrdt_update_cnt
		.p3_tx_st_hcrdt_init_ack_o   (p3_tx_st_hcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Hcrdtt_init_ack
		.p3_tx_st_dcrdt_init_i       (p3_tx_st_dcrdt_init_i),       //   input,    width = 3,                  .tx_st_Dcrdt_init
		.p3_tx_st_dcrdt_update_i     (p3_tx_st_dcrdt_update_i),     //   input,    width = 3,                  .tx_st_Dcrdt_update
		.p3_tx_st_dcrdt_update_cnt_i (p3_tx_st_dcrdt_update_cnt_i), //   input,   width = 12,                  .tx_st_Dcrdt_update_cnt
		.p3_tx_st_dcrdt_init_ack_o   (p3_tx_st_dcrdt_init_ack_o),   //  output,    width = 3,                  .tx_st_Dcrdt_init_ack
		.p3_tx_st0_hdr_o             (p3_tx_st0_hdr_o),             //  output,  width = 128,                  .tx_st0_hdr
		.p3_tx_st0_prefix_o          (p3_tx_st0_prefix_o),          //  output,   width = 32,                  .tx_st0_prefix
		.p3_tx_st0_hvalid_o          (p3_tx_st0_hvalid_o),          //  output,    width = 1,                  .tx_st0_hvalid
		.p3_tx_st0_pvalid_o          (p3_tx_st0_pvalid_o),          //  output,    width = 1,                  .tx_st0_pvalid
		.p3_tx_st1_hdr_o             (p3_tx_st1_hdr_o),             //  output,  width = 128,                  .tx_st1_hdr
		.p3_tx_st1_prefix_o          (p3_tx_st1_prefix_o),          //  output,   width = 32,                  .tx_st1_prefix
		.p3_tx_st1_hvalid_o          (p3_tx_st1_hvalid_o),          //  output,    width = 1,                  .tx_st1_hvalid
		.p3_tx_st1_pvalid_o          (p3_tx_st1_pvalid_o),          //  output,    width = 1,                  .tx_st1_pvalid
		.p0_tx_st0_ready_i           (p0_tx_st0_ready_i),           //   input,    width = 1,         p0_tx_st0.ready
		.p0_tx_st0_data_o            (p0_tx_st0_data_o),            //  output,  width = 128,                  .data
		.p0_tx_st0_sop_o             (p0_tx_st0_sop_o),             //  output,    width = 1,                  .startofpacket
		.p0_tx_st0_eop_o             (p0_tx_st0_eop_o),             //  output,    width = 1,                  .endofpacket
		.p0_tx_st0_dvalid_o          (p0_tx_st0_dvalid_o),          //  output,    width = 1,                  .valid
		.p1_tx_st0_ready_i           (p1_tx_st0_ready_i),           //   input,    width = 1,         p1_tx_st0.ready
		.p1_tx_st0_data_o            (p1_tx_st0_data_o),            //  output,  width = 128,                  .data
		.p1_tx_st0_sop_o             (p1_tx_st0_sop_o),             //  output,    width = 1,                  .startofpacket
		.p1_tx_st0_eop_o             (p1_tx_st0_eop_o),             //  output,    width = 1,                  .endofpacket
		.p1_tx_st0_dvalid_o          (p1_tx_st0_dvalid_o),          //  output,    width = 1,                  .valid
		.p2_tx_st0_ready_i           (p2_tx_st0_ready_i),           //   input,    width = 1,         p2_tx_st0.ready
		.p2_tx_st0_data_o            (p2_tx_st0_data_o),            //  output,  width = 128,                  .data
		.p2_tx_st0_sop_o             (p2_tx_st0_sop_o),             //  output,    width = 1,                  .startofpacket
		.p2_tx_st0_eop_o             (p2_tx_st0_eop_o),             //  output,    width = 1,                  .endofpacket
		.p2_tx_st0_dvalid_o          (p2_tx_st0_dvalid_o),          //  output,    width = 1,                  .valid
		.p3_tx_st0_ready_i           (p3_tx_st0_ready_i),           //   input,    width = 1,         p3_tx_st0.ready
		.p3_tx_st0_data_o            (p3_tx_st0_data_o),            //  output,  width = 128,                  .data
		.p3_tx_st0_sop_o             (p3_tx_st0_sop_o),             //  output,    width = 1,                  .startofpacket
		.p3_tx_st0_eop_o             (p3_tx_st0_eop_o),             //  output,    width = 1,                  .endofpacket
		.p3_tx_st0_dvalid_o          (p3_tx_st0_dvalid_o),          //  output,    width = 1,                  .valid
		.p0_tx_st1_data_o            (p0_tx_st1_data_o),            //  output,  width = 128,         p0_tx_st1.data
		.p0_tx_st1_sop_o             (p0_tx_st1_sop_o),             //  output,    width = 1,                  .startofpacket
		.p0_tx_st1_eop_o             (p0_tx_st1_eop_o),             //  output,    width = 1,                  .endofpacket
		.p0_tx_st1_dvalid_o          (p0_tx_st1_dvalid_o),          //  output,    width = 1,                  .valid
		.p1_tx_st1_data_o            (p1_tx_st1_data_o),            //  output,  width = 128,         p1_tx_st1.data
		.p1_tx_st1_sop_o             (p1_tx_st1_sop_o),             //  output,    width = 1,                  .startofpacket
		.p1_tx_st1_eop_o             (p1_tx_st1_eop_o),             //  output,    width = 1,                  .endofpacket
		.p1_tx_st1_dvalid_o          (p1_tx_st1_dvalid_o),          //  output,    width = 1,                  .valid
		.p2_tx_st1_data_o            (p2_tx_st1_data_o),            //  output,  width = 128,         p2_tx_st1.data
		.p2_tx_st1_sop_o             (p2_tx_st1_sop_o),             //  output,    width = 1,                  .startofpacket
		.p2_tx_st1_eop_o             (p2_tx_st1_eop_o),             //  output,    width = 1,                  .endofpacket
		.p2_tx_st1_dvalid_o          (p2_tx_st1_dvalid_o),          //  output,    width = 1,                  .valid
		.p3_tx_st1_data_o            (p3_tx_st1_data_o),            //  output,  width = 128,         p3_tx_st1.data
		.p3_tx_st1_sop_o             (p3_tx_st1_sop_o),             //  output,    width = 1,                  .startofpacket
		.p3_tx_st1_eop_o             (p3_tx_st1_eop_o),             //  output,    width = 1,                  .endofpacket
		.p3_tx_st1_dvalid_o          (p3_tx_st1_dvalid_o),          //  output,    width = 1,                  .valid
    // CSR <-> Trace Recorder
    .trace_valid_0            ( trace_valid_0 ), // Output from CSR Top
    .trace_valid_1            ( trace_valid_1 ), // Output from CSR Top
    .trace_data_0            ( trace_data_0 ), // Output from CSR Top
    .trace_data_1            ( trace_data_1 ), // Output from CSR Top
    .trace_buffer_base_addr_0            ( trace_buffer_base_addr_0 ), // Output from CSR Top
    .trace_buffer_base_addr_1            ( trace_buffer_base_addr_1 ), // Output from CSR Top
    .trace_buffer_size_0                 ( trace_buffer_size_0      ), // Output from CSR Top
    .trace_buffer_size_1                 ( trace_buffer_size_1      ), // Output from CSR Top
    .control_register_0                  ( control_register_0       ), // Output from CSR Top
    .control_register_1                  ( control_register_1       ), // Output from CSR Top
    .dropped_traces_0                    ( dropped_traces_0         ), // Input to CSR Top
    .dropped_traces_1                    ( dropped_traces_1         ), // Input to CSR Top
    .written_traces_0                    ( written_traces_0         ), // Input to CSR Top
    .written_traces_1                    ( written_traces_1         )  // Input to CSR Top
	);

endmodule
